// Jacob Panov
// lab01_data yapp UVC package for accelerated UVM
// yapp_pkg.sv

package yapp_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "/home/jpanov/Cadence/uvma_training_1.2.6rev1/uvm/lab01_data/sv/yapp_packet.sv"

    
endpackage : yapp_pkg