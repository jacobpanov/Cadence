// Jacob Panov
// lab01_data yapp UVC package for accelerated UVM
// yapp_pkg.sv

package yapp_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "yapp_packet.sv"
  
endpackage